library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity regPC is
	port
	(
		ck,rst: in std_logic;
		pc : in std_logic_vector(31 downto 0);
		
	);
end regPC;

architecture Behavioral of regPC is

begin


end Behavioral;

